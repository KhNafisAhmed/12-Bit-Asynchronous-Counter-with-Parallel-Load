class bc_tr_item;
  
  //Inputs
  logic enable;
  logic reset_n;
  logic load;
  logic up_down;
  logic [11:0]data;
  
  //Outputs
  logic [11:0]count;
  
endclass