`include "COUNTER_12bit.sv"
`include "bc_tr_item.sv"
`include "bc_driver.sv"
`include "bc_monitor.sv"
`include "bc_scb.sv"
`include "bc_agent.sv"
`include "bc_env.sv"
`include "bc_test.sv"
`include "bc_interface.sv"